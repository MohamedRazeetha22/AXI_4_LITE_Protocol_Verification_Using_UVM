`ifndef AXI_ENVIRONMENT
`define AXI_ENVIRONMENT
class axi_environment extends uvm_env;
`uvm_component_utils (axi_environment)
axi_agent agt;
axi_scoreboard scb;
// axi_coverage cov;
function new (string name="axi_environment", uvm_component parent);
super.new(name, parent);
endfunction
function void build_phase (uvm_phase phase);
super.build_phase (phase);
agt=axi_agent::type_id::create("agt",this);
scb=axi_scoreboard::type_id::create("scb",this);
// cov=axi_coverage:: type_id::create("cov",this);
endfunction
function void connect_phase (uvm_phase phase);
agt.mon.ap.connect(scb.analysis_export);
// agt.mon.ap.connect(cov.analysis_export);
endfunction
endclass
`endif
