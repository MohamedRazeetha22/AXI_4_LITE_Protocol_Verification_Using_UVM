`ifndef AXI_ENVIRONMENT_PKG
`define AXI_ENVIRONMENT_PKG
package axi_environment_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
import axi_agent_pkg::*;
`include "axi_scoreboard.sv"
//`include "axi_coverage.sv"
`include "axi_environment.sv"
endpackage
`endif
